`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/03/28 19:36:42
// Design Name: 
// Module Name: tb_phase_a_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_phase_a#(
    parameter M_SIZE = 3072,
    parameter RADIX = 72,
    parameter SIZE_LOG = 6,
    parameter FIFO_DEPTH = 4,
    parameter FIFO_AddrWidth = 3,
    parameter SIZE_ADD = 128*25
)(
    );
    reg clk, rst_n, en;
    reg [3149:0] a;
    reg [3071:0] m;
    reg [3073:0] m_n;
    reg [79:0] m_prime;
    reg if_last;
    wire [3071:0] new_a;
    wire [2:0] cnt_4;
    wire en_out;
    
    initial begin
        clk = 0;
        rst_n = 0;
        en = 0;
        a = 3144'h5537b809d650de8821a83a5433a9d61aede0b5920116118d86fb93a8d61ff5a55a3e1a86a9120ba88af0ff4819be8672a58ecbc4400842af1066a7b2e35e526d9ab97bd64db7bff40899184841441aa17a2d7841cf20bc9a5fc943298506d301af280f381f7926c35def357682db8c4db8efe60f0aa935118ab780d2973963903eb6d14bb6540990f80c8061362db2be2bf1cc084dce716c58cca95c5cd0c1b936019cd4759e88ad73f4da76a03fbeef68cb9e02460732361921f86cce6536ba073754de30ed0e06ed36943c5ec050f7ddd4257fbb5af45a6f419c93f11cd49134357a0be4edc9ec3ca2f8b87afa9fa492ab0d79195a0fee32d288531fef019fa0c99c50fed25f253cb31035ef94ecbf2d1565bdc8cc519313cbef7757b04f50f8ca834effd0688af300f3659a9447316b59e67540d31c8be01cb54ecae0e8ca60cf668014db967669e48796ecd0807113b29d0a42eb574f2e554879c44eb5d200585ffbd15b31f5f7a0a3a557a31bc8400bf88f4748907725c7be2d13da5531000000000000000000;
        m = 3072'hdc85279b3f9f6f56ed70ec798632ff7f62829f9aed27ce9b97bf748a8768c48364a1f91bacfdd03d5190b29661de1d3d206b56c498e67cafbee993abecc98f843cdc450214c40389a03b958e0fcceeacdc05af7438ba1a595c3e7931966a71299fbaedda383a619433cc35a51da18d6acc030a84b25333a327328ca85b44e416ccb17ae7676587791240ca9c49d1cf8218a83e6560bd24eeca83e1bae2e7ea0d8f7ad7f578fb28cc66ea66547c8b99954ca77217d79e0d40cf15e92a1da2bc22c1ff04bab3064e192857ae677f43bf3f1e52b96d702283a7dc9988476fa7ad499f015f0dd2b5d4422762d34c42635dbc83c14fdedef8f76bbe1ad03d2c60075887f5811f7765d9ae7d4201524cd355e8d8e73925526c356eb8f676af0217a64b74cb4ad6525fc9f7fca40ef0ee70f11022804bd7bf7c2321c9505c6ab348082a84955d0a38f8dda6e8c347268de733f4adf6475bf4dbf88443f43365070d2d21c472527036376a0baf155d8bf192f20254882416f304ad08992cc4e36483d004;
        m_n = 3074'h3237ad864c06090a9128f138679cd00809d7d606512d8316468408b7578973b7c9b5e06e453022fc2ae6f4d699e21e2c2df94a93b6719835041166c541336707bc323bafdeb3bfc765fc46a71f033115323fa508bc745e5a6a3c186ce69958ed660451225c7c59e6bcc33ca5ae25e729533fcf57b4daccc5cd8cd7357a4bb1be9334e8518989a7886edbf3563b62e307de757c19a9f42db11357c1e451d1815f27085280a8704d733991599ab8374666ab3588de82861f2bf30ea16d5e25d43dd3e00fb454cf9b1e6d7a8519880bc40c0e1ad46928fdd7c58236677b8905852b660fea0f22d4a2bbdd89d2cb3bd9ca2437c3eb0212107089441e52fc2d39ff8a7780a7ee0889a265182bdfeadb32caa172718c6daad93ca9147098950fde859b48b34b529ada03608035bf10f118f0eefdd7fb4284083dcde36afa3954cb7f7d57b6aa2f5c7072259173cb8d97218cc0b5209b8a40b24077bbc0bcc9af8f2d2de3b8dad8fc9c895f450eaa2740e6d0dfdab77dbe90cfb52f766d33b1c9b7c2ffc;
        m_prime = 80'h4a4c0ccb4cb4e139f56b;
        if_last = 1;
        #15
        a=a<<6;
        rst_n = 1;
        #20
        en = 1;
        // time 195 ns
        // answer 3072'hd0a359e4d59ad93c86094ea7fc4baa9b2c3a54ee0599a193484ef2e2ddfa992d14c4b0e6a44cc6e817d1d8ed943053b6271e948a06e264af804c0cfdf516fd6cd7f4b8c8609c25406e23a9d69bd7e00f727284fa5b1ad185d1b98326205de202099f4235a6d048c73837803acb5ab733a53b94076fa0def1c3e427971658df7c12046426d4560a68dd022d723c58041ae769f7727778ccc813b6edd0cb24f3a7c13ac1fd9548c4b536a17d461cc1ba441e163c6af7bccc0a848d074e9fe313ce9e7b2c4775a9b8c9e34f6c4a74f7e318fab487e2711fa31e389a8e186d8fb34976546ce3c365253f0d039d5e4514f9dc080c993e8ab72fb51482d2a89919efa56f946e34d2452d370f6d64d1e5309df1fdd6bab1ec117083ba0a52cfc836896b6375799eb7803bf6b23373e72f58322722fd15529285015137fa3004fb3e36957bdb146094a504799aafbc89756d5dcd4e6587ec8967af18f6450a354da97914a8b9b757d8971afbd1d9713044ec0f7e71b096a9fe6a4eb67a8f5c8ef7358ba0
        #10;
        en = 0;
        #30
        a = 3144'h5547b809d650de8821a83a5433a9d61aede0b5920116118d86fb93a8d61ff5a55a3e1a86a9120ba88af0ff4819be8672a58ecbc4400842af1066a7b2e35e526d9ab97bd64db7bff40899184841441aa17a2d7841cf20bc9a5fc943298506d301af280f381f7926c35def357682db8c4db8efe60f0aa935118ab780d2973963903eb6d14bb6540990f80c8061362db2be2bf1cc084dce716c58cca95c5cd0c1b936019cd4759e88ad73f4da76a03fbeef68cb9e02460732361921f86cce6536ba073754de30ed0e06ed36943c5ec050f7ddd4257fbb5af45a6f419c93f11cd49134357a0be4edc9ec3ca2f8b87afa9fa492ab0d79195a0fee32d288531fef019fa0c99c50fed25f253cb31035ef94ecbf2d1565bdc8cc519313cbef7757b04f50f8ca834effd0688af300f3659a9447316b59e67540d31c8be01cb54ecae0e8ca60cf668014db967669e48796ecd0807113b29d0a42eb574f2e554879c44eb5d200585ffbd15b31f5f7a0a3a557a31bc8400bf88f4748907725c7be2d13da5531000000000000000000;
        en = 1;
        // time 235 ns
        // answer 3072'hc1efd103483c33684a0016b5ef3ba62e7e021a82bf725c121cf5f7eaefb03c6da2cfda13dbf575ecf89a5deef0db57dd99aefa2831f97610677a68cdbdecd51fa7e33bbaca7720cbb064304f98160983798b1fb163d1d15a1f61ed7091333ec74b127b2a8a67cad3520562a355c1531be241db63f05f0a3243282d97d3b83f9246f5c8b6693b803db21276508e8224b441aa15e9c9df26f904e7b90e6dc69c0476264510053e951d93f445fd1db4f2e73a8830880b510cd5b5a158bbf436006f00afbaf168bf3d783fe0cff5acee5f4338ad191733b7ec7a5532e71eb474a27b1668252562e8f98ef77fb83ab81d8c7bd97291a98a4021a42f528429ff9e40de3e4b189319ee29b670c90c6bf971a865ca838a38dedb99f9b89d8eb2675c4b857e3bfeb01d3ce90b53d0f6bef870eb8586d747c5d81199b04b3def1e708846dd5fa014bbb218e6d71b68221cafe3679f583a7556018509ecbdcebe40fc943faf30f1046789a8ede9796f4ee8949848ef921e39453460e1efad594f9b2f3002f8
        if_last = 0;
        #10 en = 0;
        #1000; 
        $finish;
    end


    always #5 clk = ~clk;
    phase_a #(
    .Size(M_SIZE), 
    .radix(RADIX), 
    .Size_log(SIZE_LOG), 
    .Size_add(SIZE_ADD))
    phase_a(.clk(clk), .rst_n(rst_n), .a(a), .m(m), .m_n(m_n), .m_prime(m_prime), .en(en), .if_last(if_last), .new_a(new_a), .cnt_4(cnt_4), .en_out(en_out));
endmodule
